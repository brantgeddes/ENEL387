** Profile: "SCHEMATIC1-387ZFC_Sim"  [ C:\Users\brant\Desktop\School\Sem 7\ENEL 387\Project\Sims\387ZFC_Sim-PSpiceFiles\SCHEMATIC1\387ZFC_Sim.sim ] 

** Creating circuit file "387ZFC_Sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\brant\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 100mS 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
